(* Compatibility of Require with backtracking at interactive module end *)

Module A.
Require ListDef.
End A.
