(* Compatibility of Require with backtracking at interactive module end *)

Module A.
Require List.
End A.
